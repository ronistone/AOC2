library IEEE; 
use IEEE.STD_LOGIC_1164.all;

entity exercise1 is
	port(	a, b, c: in STD_LOGIC;
			y, z: out STD_LOGIC);
end;

architecture synth of exercise1 is
begin
	y <= (a and b and c) or (a and b and not c) or (a and not b and c);
	z <= (a and b) or (not a and not b);
end;